`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:12:30 05/15/2016 
// Design Name: 
// Module Name:    IM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module IM(IAddr,
			InsMemRW,
			DataOut
			);
	input[31:0] IAddr;
	input InsMemRW;
	
	output reg[31:0] DataOut;
	
	reg[7:0] rom[0:255];
	
	initial
		begin
			// j   0x0000 0064
			rom[32'h00000028] <= 8'b11100000;
			rom[32'h00000029] <= 8'b00000000;
			rom[32'h0000002a] <= 8'b00000000;
			rom[32'h0000002b] <= 8'b00011001;
			// ori  $1, $0, 8
			rom[32'h00000064] <= 8'b01001000;
			rom[32'h00000065] <= 8'b00000001;
			rom[32'h00000066] <= 8'b00000000;
			rom[32'h00000067] <= 8'b00001000;
			// addi $2, $0, 7
			rom[32'h00000068] <= 8'b00001000;
			rom[32'h00000069] <= 8'b00000010;
			rom[32'h0000006a] <= 8'b00000000;
			rom[32'h0000006b] <= 8'b00000111;
			// sub $3, $1, $2
			rom[32'h0000006c] <= 8'b00000100;
			rom[32'h0000006d] <= 8'b00100010;
			rom[32'h0000006e] <= 8'b00011000;
			rom[32'h0000006f] <= 8'b00000000;
			// add $4, $1, $2
			rom[32'h00000070] <= 8'b00000000;
			rom[32'h00000071] <= 8'b00100010;
			rom[32'h00000072] <= 8'b00100000;
			rom[32'h00000073] <= 8'b00000000;
			// and $5, $2, $4
			rom[32'h00000074] <= 8'b01000100;
			rom[32'h00000075] <= 8'b01000100;
			rom[32'h00000076] <= 8'b00101000;
			rom[32'h00000077] <= 8'b00000000;
			// or $6, $1, $3
			rom[32'h00000078] <= 8'b01000000;
			rom[32'h00000079] <= 8'b00100011;
			rom[32'h0000007a] <= 8'b00110000;
			rom[32'h0000007b] <= 8'b00000000;
			// move $7, $1
			rom[32'h0000007c] <= 8'b10000000;
			rom[32'h0000007d] <= 8'b00100000;
			rom[32'h0000007e] <= 8'b00111000;
			rom[32'h0000007f] <= 8'b00000000;
			// jal  0x0000 0098
			rom[32'h00000080] <= 8'b11101000;
			rom[32'h00000081] <= 8'b00000000;
			rom[32'h00000082] <= 8'b00000000;
			rom[32'h00000083] <= 8'b00100110;
			// slt $8, $1, $2
			rom[32'h00000084] <= 8'b10011100;
			rom[32'h00000085] <= 8'b00100010;
			rom[32'h00000086] <= 8'b01000000;
			rom[32'h00000087] <= 8'b00000000;
			// slt $9, $1, $4
			rom[32'h00000088] <= 8'b10011100;
			rom[32'h00000089] <= 8'b00100100;
			rom[32'h0000008a] <= 8'b01001000;
			rom[32'h0000008b] <= 8'b00000000;
			// sll $3, $3, 3
			rom[32'h0000008c] <= 8'b01100000;
			rom[32'h0000008d] <= 8'b01100000;
			rom[32'h0000008e] <= 8'b00011000;
			rom[32'h0000008f] <= 8'b11000000;
			// beq $3, $1, -2 ת8C
			rom[32'h00000090] <= 8'b11010000;
			rom[32'h00000091] <= 8'b01100001;
			rom[32'h00000092] <= 8'b11111111;
			rom[32'h00000093] <= 8'b11111110;
			// halt
			rom[32'h00000094] <= 8'b11111100;
			rom[32'h00000095] <= 8'b00000000;
			rom[32'h00000096] <= 8'b00000000;
			rom[32'h00000097] <= 8'b00000000;
			// sw $6, 1($2)
			rom[32'h00000098] <= 8'b11000000;
			rom[32'h00000099] <= 8'b01000110;
			rom[32'h0000009a] <= 8'b00000000;
			rom[32'h0000009b] <= 8'b00000001;
			// lw $11, 1($2)
			rom[32'h0000009c] <= 8'b11000100;
			rom[32'h0000009d] <= 8'b01001011;
			rom[32'h0000009e] <= 8'b00000000;
			rom[32'h0000009f] <= 8'b00000001;
			// jr  $31
			rom[32'h000000a0] <= 8'b11100111;
			rom[32'h000000a1] <= 8'b11100000;
			rom[32'h000000a2] <= 8'b00000000;
			rom[32'h000000a3] <= 8'b00000000;
		end
	
	always @(InsMemRW or IAddr)
		begin
			if (InsMemRW == 0)
				DataOut = {rom[IAddr][7:0], rom[IAddr + 1][7:0], rom[IAddr + 2][7:0], rom[IAddr + 3][7:0]};
		end	
endmodule














